package globals;
  parameter int DW=8;
  parameter int CW=4;
endpackage
